`timescale 1ns/1ps
module c880_test (gat1, gat8, gat13, gat17, gat26, gat29, gat36, gat42, gat51, gat55, gat59, gat68, gat72, gat73, gat74, gat75, gat80, gat85, gat86, gat87, gat88, gat89, gat90, gat91, gat96, gat101, gat106, gat111, gat116, gat121, gat126, gat130, gat135, gat138, gat143, gat146, gat149, gat152, gat153, gat156, gat159, gat165, gat171, gat177, gat183, gat189, gat195, gat201, gat207, gat210, gat219, gat228, gat237, gat246, gat255, gat259, gat260, gat261, gat267, gat268, input gat1, gat8, gat13, gat17, gat26, gat29, gat36, gat42, gat51, gat55, gat59, gat68, gat72, gat73, gat74, gat75, gat80, gat85, gat86, gat87, gat88, gat89, gat90, gat91, gat96, gat101, gat106, gat111, gat116, gat121, gat126, gat130, gat135, gat138, gat143, gat146, gat149, gat152, gat153, gat156, gat159, gat165, gat171, gat177, gat183, gat189, gat195, gat201, gat207, gat210, gat219, gat228, gat237, gat246, gat255, gat259, gat260, gat261, gat267, gat268;
output wire gat2, gat3, gat4, gat5, gat6, gat7, gat9, gat10, gat11, gat12, gat14, gat15, gat16, gat18, gat19, gat20, gat21, gat22, gat23, gat24, gat25, gat27, gat28, gat30, gat31, gat32, gat33, gat34, gat35, gat37, gat38, gat39, gat40, gat41, gat43, gat44, gat45, gat46, gat47, gat48, gat49, gat50, gat52, gat53, gat54, gat56, gat57, gat58, gat60, gat61, gat62, gat63, gat64, gat65, gat66, gat67, gat69, gat70, gat71, gat76, gat77, gat78, gat79, gat81, gat82, gat83, gat84, gat92, gat93, gat94, gat95, gat97, gat98, gat99, gat100, gat102, gat103, gat104, gat105, gat107, gat108, gat109, gat110, gat112, gat113, gat114, gat115, gat117, gat118, gat119, gat120, gat122, gat123, gat124, gat125, gat127, gat128, gat129, gat131, gat132, gat133, gat134, gat136, gat137, gat139, gat140, gat141, gat142, gat144, gat145, gat147, gat148, gat150, gat151, gat154, gat155, gat157, gat158, gat160, gat161, gat162, gat163, gat164, gat166, gat167, gat168, gat169, gat170, gat172, gat173, gat174, gat175, gat176, gat178, gat179, gat180, gat181, gat182, gat184, gat185, gat186, gat187, gat188, gat190, gat191, gat192, gat193, gat194, gat196, gat197, gat198, gat199, gat200, gat202, gat203, gat204, gat205, gat206, gat208, gat209, gat211, gat212, gat213, gat214, gat215, gat216, gat217, gat218, gat220, gat221, gat222, gat223, gat224, gat225, gat226, gat227, gat229, gat230, gat231, gat232, gat233, gat234, gat235, gat236, gat238, gat239, gat240, gat241, gat242, gat243, gat244, gat245, gat247, gat248, gat249, gat250, gat251, gat252, gat253, gat254, gat256, gat257, gat258, gat262, gat263, gat264, gat265, gat266, gat269, gat270, gat271, gat272, gat273, gat274, gat275, gat276, gat277, gat278, gat279, gat280, gat281, gat282, gat283, gat284, gat285, gat286, gat287, gat288, gat289, gat290, gat291, gat292, gat293, gat294, gat295, gat296, gat297, gat298, gat299, gat300, gat301, gat302, gat303, gat304, gat305, gat306, gat307, gat308, gat309, gat310, gat311, gat312, gat313, gat314, gat315, gat316, gat317, gat318, gat319, gat320, gat321, gat322, gat323, gat324, gat325, gat326, gat327, gat328, gat329, gat330, gat331, gat332, gat333, gat334, gat335, gat336, gat337, gat338, gat339, gat340, gat341, gat342, gat343, gat344, gat345, gat346, gat347, gat348, gat349, gat350, gat351, gat352, gat353, gat354, gat355, gat356, gat357, gat358, gat359, gat360, gat361, gat362, gat363, gat364, gat365, gat366, gat367, gat368, gat369, gat370, gat371, gat372, gat373, gat374, gat375, gat376, gat377, gat378, gat379, gat380, gat381, gat382, gat383, gat384, gat385, gat386, gat387, gat392, gat393, gat394, gat395, gat396, gat397, gat398, gat399, gat400, gat401, gat402, gat403, gat404, gat405, gat406, gat407, gat408, gat409, gat410, gat411, gat412, gat413, gat414, gat415, gat416, gat417, gat424, gat425, gat426, gat427, gat428, gat429, gat430, gat431, gat432, gat433, gat434, gat435, gat436, gat437, gat438, gat439, gat440, gat441, gat442, gat443, gat444, gat445, gat451, gat452, gat453, gat454, gat455, gat456, gat457, gat458, gat459, gat460, gat461, gat462, gat463, gat464, gat465, gat466, gat467, gat468, gat469, gat470, gat471, gat472, gat473, gat474, gat475, gat476, gat477, gat478, gat479, gat480, gat481, gat482, gat483, gat484, gat485, gat486, gat487, gat488, gat489, gat490, gat491, gat492, gat493, gat494, gat495, gat496, gat497, gat498, gat499, gat500, gat501, gat502, gat503, gat504, gat505, gat506, gat507, gat508, gat509, gat510, gat511, gat512, gat513, gat514, gat515, gat516, gat517, gat518, gat519, gat520, gat521, gat522, gat523, gat524, gat525, gat526, gat527, gat528, gat529, gat530, gat531, gat532, gat533, gat534, gat535, gat536, gat537, gat538, gat539, gat540, gat541, gat542, gat543, gat544, gat545, gat546, gat547, gat548, gat549, gat550, gat551, gat552, gat553, gat554, gat555, gat556, gat557, gat558, gat559, gat560, gat561, gat562, gat563, gat564, gat565, gat566, gat567, gat568, gat569, gat570, gat571, gat572, gat573, gat574, gat575, gat576, gat577, gat578, gat579, gat580, gat581, gat582, gat583, gat584, gat585, gat586, gat587, gat588, gat589, gat590, gat591, gat592, gat593, gat594, gat595, gat596, gat597, gat598, gat599, gat600, gat601, gat602, gat603, gat604, gat605, gat606, gat607, gat608, gat609, gat610, gat611, gat612, gat613, gat614, gat615, gat616, gat617, gat618, gat619, gat620, gat621, gat622, gat623, gat624, gat625, gat626, gat627, gat628, gat629, gat630, gat631, gat632, gat633, gat634, gat635, gat636, gat637, gat638, gat639, gat640, gat641, gat642, gat643, gat644, gat645, gat646, gat647, gat648, gat649, gat650, gat651, gat652, gat653, gat654, gat655, gat656, gat657, gat658, gat659, gat660, gat661, gat662, gat663, gat664, gat665, gat666, gat667, gat668, gat669, gat670, gat671, gat672, gat673, gat674, gat675, gat676, gat677, gat678, gat679, gat680, gat681, gat682, gat683, gat684, gat685, gat686, gat687, gat688, gat689, gat690, gat691, gat692, gat693, gat694, gat695, gat696, gat697, gat698, gat699, gat700, gat701, gat702, gat703, gat704, gat705, gat706, gat707, gat708, gat709, gat710, gat711, gat712, gat713, gat714, gat715, gat716, gat717, gat718, gat719, gat720, gat721, gat722, gat723, gat724, gat725, gat726, gat727, gat728, gat729, gat730, gat731, gat732, gat733, gat734, gat735, gat736, gat737, gat738, gat739, gat740, gat741, gat742, gat743, gat744, gat745, gat746, gat747, gat748, gat749, gat750, gat751, gat752, gat753, gat754, gat755, gat756, gat757, gat758, gat759, gat760, gat761, gat762, gat763, gat764, gat765, gat766, gat769, gat770, gat771, gat772, gat773, gat774, gat775, gat776, gat777, gat778, gat779, gat780, gat781, gat782, gat783, gat784, gat785, gat786, gat787, gat788, gat789, gat790, gat791, gat792, gat793, gat794, gat795, gat796, gat797, gat798, gat799, gat800, gat801, gat802, gat803, gat804, gat805, gat806, gat807, gat808, gat809, gat810, gat811, gat812, gat813, gat814, gat815, gat816, gat817, gat818, gat819, gat820, gat821, gat822, gat823, gat824, gat825, gat826, gat827, gat828, gat829, gat830, gat831, gat832, gat833, gat834, gat835, gat836, gat837, gat838, gat839, gat840, gat841, gat842, gat843, gat844, gat845, gat846, gat847, gat848, gat849, gat851, gat852, gat853, gat854, gat855, gat856, gat857, gat858, gat859, gat860, gat861, gat862, gat867, gat868, gat869, gat870, gat871, gat872, gat873, gat875, gat876, gat877;
assign gat2 = gat1;
assign gat3 = gat1;
assign gat4 = gat1;
assign gat5 = gat1;
assign gat6 = gat1;
assign gat7 = gat1;
assign gat9 = gat8;
assign gat10 = gat8;
assign gat11 = gat8;
assign gat12 = gat8;
assign gat14 = gat13;
assign gat15 = gat13;
assign gat16 = gat13;
assign gat18 = gat17;
assign gat19 = gat17;
assign gat20 = gat17;
assign gat21 = gat17;
assign gat22 = gat17;
assign gat23 = gat17;
assign gat24 = gat17;
assign gat25 = gat17;
assign gat27 = gat26;
assign gat28 = gat26;
assign gat30 = gat29;
assign gat31 = gat29;
assign gat32 = gat29;
assign gat33 = gat29;
assign gat34 = gat29;
assign gat35 = gat29;
assign gat37 = gat36;
assign gat38 = gat36;
assign gat39 = gat36;
assign gat40 = gat36;
assign gat41 = gat36;
assign gat43 = gat42;
assign gat44 = gat42;
assign gat45 = gat42;
assign gat46 = gat42;
assign gat47 = gat42;
assign gat48 = gat42;
assign gat49 = gat42;
assign gat50 = gat42;
assign gat52 = gat51;
assign gat53 = gat51;
assign gat54 = gat51;
assign gat56 = gat55;
assign gat57 = gat55;
assign gat58 = gat55;
assign gat60 = gat59;
assign gat61 = gat59;
assign gat62 = gat59;
assign gat63 = gat59;
assign gat64 = gat59;
assign gat65 = gat59;
assign gat66 = gat59;
assign gat67 = gat59;
assign gat69 = gat68;
assign gat70 = gat68;
assign gat71 = gat68;
assign gat76 = gat75;
assign gat77 = gat75;
assign gat78 = gat75;
assign gat79 = gat75;
assign gat81 = gat80;
assign gat82 = gat80;
assign gat83 = gat80;
assign gat84 = gat80;
assign gat92 = gat91;
assign gat93 = gat91;
assign gat94 = gat91;
assign gat95 = gat91;
assign gat97 = gat96;
assign gat98 = gat96;
assign gat99 = gat96;
assign gat100 = gat96;
assign gat102 = gat101;
assign gat103 = gat101;
assign gat104 = gat101;
assign gat105 = gat101;
assign gat107 = gat106;
assign gat108 = gat106;
assign gat109 = gat106;
assign gat110 = gat106;
assign gat112 = gat111;
assign gat113 = gat111;
assign gat114 = gat111;
assign gat115 = gat111;
assign gat117 = gat116;
assign gat118 = gat116;
assign gat119 = gat116;
assign gat120 = gat116;
assign gat122 = gat121;
assign gat123 = gat121;
assign gat124 = gat121;
assign gat125 = gat121;
assign gat127 = gat126;
assign gat128 = gat126;
assign gat129 = gat126;
assign gat131 = gat130;
assign gat132 = gat130;
assign gat133 = gat130;
assign gat134 = gat130;
assign gat136 = gat135;
assign gat137 = gat135;
assign gat139 = gat138;
assign gat140 = gat138;
assign gat141 = gat138;
assign gat142 = gat138;
assign gat144 = gat143;
assign gat145 = gat143;
assign gat147 = gat146;
assign gat148 = gat146;
assign gat150 = gat149;
assign gat151 = gat149;
assign gat154 = gat153;
assign gat155 = gat153;
assign gat157 = gat156;
assign gat158 = gat156;
assign gat160 = gat159;
assign gat161 = gat159;
assign gat162 = gat159;
assign gat163 = gat159;
assign gat164 = gat159;
assign gat166 = gat165;
assign gat167 = gat165;
assign gat168 = gat165;
assign gat169 = gat165;
assign gat170 = gat165;
assign gat172 = gat171;
assign gat173 = gat171;
assign gat174 = gat171;
assign gat175 = gat171;
assign gat176 = gat171;
assign gat178 = gat177;
assign gat179 = gat177;
assign gat180 = gat177;
assign gat181 = gat177;
assign gat182 = gat177;
assign gat184 = gat183;
assign gat185 = gat183;
assign gat186 = gat183;
assign gat187 = gat183;
assign gat188 = gat183;
assign gat190 = gat189;
assign gat191 = gat189;
assign gat192 = gat189;
assign gat193 = gat189;
assign gat194 = gat189;
assign gat196 = gat195;
assign gat197 = gat195;
assign gat198 = gat195;
assign gat199 = gat195;
assign gat200 = gat195;
assign gat202 = gat201;
assign gat203 = gat201;
assign gat204 = gat201;
assign gat205 = gat201;
assign gat206 = gat201;
assign gat208 = gat207;
assign gat209 = gat207;
assign gat211 = gat210;
assign gat212 = gat210;
assign gat213 = gat210;
assign gat214 = gat210;
assign gat215 = gat210;
assign gat216 = gat210;
assign gat217 = gat210;
assign gat218 = gat210;
assign gat220 = gat219;
assign gat221 = gat219;
assign gat222 = gat219;
assign gat223 = gat219;
assign gat224 = gat219;
assign gat225 = gat219;
assign gat226 = gat219;
assign gat227 = gat219;
assign gat229 = gat228;
assign gat230 = gat228;
assign gat231 = gat228;
assign gat232 = gat228;
assign gat233 = gat228;
assign gat234 = gat228;
assign gat235 = gat228;
assign gat236 = gat228;
assign gat238 = gat237;
assign gat239 = gat237;
assign gat240 = gat237;
assign gat241 = gat237;
assign gat242 = gat237;
assign gat243 = gat237;
assign gat244 = gat237;
assign gat245 = gat237;
assign gat247 = gat246;
assign gat248 = gat246;
assign gat249 = gat246;
assign gat250 = gat246;
assign gat251 = gat246;
assign gat252 = gat246;
assign gat253 = gat246;
assign gat254 = gat246;
assign gat256 = gat255;
assign gat257 = gat255;
assign gat258 = gat255;
assign gat262 = gat261;
assign gat263 = gat261;
assign gat264 = gat261;
assign gat265 = gat261;
assign gat266 = gat261;
nand 269gat (gat269, gat2, gat9, gat14, gat18);
nand 270gat (gat270, gat3, gat27, gat15, gat19);
assign gat271 = gat270;
assign gat272 = gat270;
and 273gat (gat273, gat30, gat37, gat43);
assign gat274 = gat273;
assign gat275 = gat273;
and 276gat (gat276, gat4, gat28, gat52);
assign gat277 = gat276;
assign gat278 = gat276;
nand 279gat (gat279, gat5, gat10, gat53, gat20);
nand 280gat (gat280, gat6, gat11, gat16, gat56);
assign gat281 = gat280;
assign gat282 = gat280;
assign gat283 = gat280;
nand 284gat (gat284, gat60, gat44, gat69, gat72);
nand 285gat (gat285, gat31, gat70);
nand 286gat (gat286, gat61, gat71, gat74);
and 287gat (gat287, gat32, gat76, gat81);
assign gat288 = gat287;
assign gat289 = gat287;
and 290gat (gat290, gat33, gat77, gat45);
and 291gat (gat291, gat34, gat38, gat82);
and 292gat (gat292, gat35, gat39, gat46);
and 293gat (gat293, gat62, gat78, gat83);
and 294gat (gat294, gat63, gat79, gat47);
and 295gat (gat295, gat64, gat40, gat84);
and 296gat (gat296, gat65, gat41, gat48);
and 297gat (gat297, gat85, gat86);
or 298gat (gat298, gat87, gat88);
assign gat299 = gat298;
assign gat300 = gat298;
nand 301gat (gat301, gat92, gat97);
or 302gat (gat302, gat93, gat98);
nand 303gat (gat303, gat102, gat107);
or 304gat (gat304, gat103, gat108);
nand 305gat (gat305, gat112, gat117);
or 306gat (gat306, gat113, gat118);
nand 307gat (gat307, gat122, gat127);
or 308gat (gat308, gat123, gat128);
and 309gat (gat309, gat12, gat139);
not 310gat (gat310, gat268);
assign gat311 = gat310;
assign gat312 = gat310;
assign gat313 = gat310;
assign gat314 = gat310;
assign gat315 = gat310;
and 316gat (gat316, gat54, gat140);
and 317gat (gat317, gat21, gat141);
and 318gat (gat318, gat152, gat142);
nand 319gat (gat319, gat66, gat157);
assign gat320 = gat319;
assign gat321 = gat319;
nor 322gat (gat322, gat22, gat49);
and 323gat (gat323, gat23, gat50);
nand 324gat (gat324, gat160, gat166);
or 325gat (gat325, gat161, gat167);
nand 326gat (gat326, gat172, gat178);
or 327gat (gat327, gat173, gat179);
nand 328gat (gat328, gat184, gat190);
or 329gat (gat329, gat185, gat191);
nand 330gat (gat330, gat196, gat202);
or 331gat (gat331, gat197, gat203);
and 332gat (gat332, gat211, gat94);
and 333gat (gat333, gat212, gat99);
and 334gat (gat334, gat213, gat104);
and 335gat (gat335, gat214, gat109);
and 336gat (gat336, gat215, gat114);
and 337gat (gat337, gat256, gat259);
and 338gat (gat338, gat216, gat119);
and 339gat (gat339, gat257, gat260);
and 340gat (gat340, gat217, gat124);
and 341gat (gat341, gat258, gat267);
not 342gat (gat342, gat269);
not 343gat (gat343, gat274);
or 344gat (gat344, gat271, gat275);
not 345gat (gat345, gat277);
not 346gat (gat346, gat278);
not 347gat (gat347, gat279);
nor 348gat (gat348, gat281, gat284);
or 349gat (gat349, gat282, gat285);
or 350gat (gat350, gat283, gat286);
not 351gat (gat351, gat293);
not 352gat (gat352, gat294);
not 353gat (gat353, gat295);
not 354gat (gat354, gat296);
nand 355gat (gat355, gat89, gat299);
and 356gat (gat356, gat90, gat300);
nand 357gat (gat357, gat301, gat302);
assign gat358 = gat357;
assign gat359 = gat357;
nand 360gat (gat360, gat303, gat304);
assign gat361 = gat360;
assign gat362 = gat360;
nand 363gat (gat363, gat305, gat306);
assign gat364 = gat363;
assign gat365 = gat363;
nand 366gat (gat366, gat307, gat308);
assign gat367 = gat366;
assign gat368 = gat366;
not 369gat (gat369, gat311);
assign gat370 = gat369;
assign gat371 = gat369;
assign gat372 = gat369;
assign gat373 = gat369;
assign gat374 = gat369;
nor 375gat (gat375, gat322, gat323);
nand 376gat (gat376, gat324, gat325);
assign gat377 = gat376;
assign gat378 = gat376;
nand 379gat (gat379, gat326, gat327);
assign gat380 = gat379;
assign gat381 = gat379;
nand 382gat (gat382, gat328, gat329);
assign gat383 = gat382;
assign gat384 = gat382;
nand 385gat (gat385, gat330, gat331);
assign gat386 = gat385;
assign gat387 = gat385;
or 392gat (gat392, gat272, gat343);
not 393gat (gat393, gat345);
assign gat394 = gat393;
assign gat395 = gat393;
assign gat396 = gat393;
assign gat397 = gat393;
assign gat398 = gat393;
not 399gat (gat399, gat346);
and 400gat (gat400, gat348, gat73);
not 401gat (gat401, gat349);
not 402gat (gat402, gat350);
not 403gat (gat403, gat355);
not 404gat (gat404, gat358);
not 405gat (gat405, gat361);
and 406gat (gat406, gat359, gat362);
not 407gat (gat407, gat364);
not 408gat (gat408, gat367);
and 409gat (gat409, gat365, gat368);
nand 410gat (gat410, gat347, gat352);
not 411gat (gat411, gat377);
not 412gat (gat412, gat380);
and 413gat (gat413, gat378, gat381);
not 414gat (gat414, gat383);
not 415gat (gat415, gat386);
and 416gat (gat416, gat384, gat387);
and 417gat (gat417, gat218, gat370);
not 424gat (gat424, gat400);
and 425gat (gat425, gat404, gat405);
and 426gat (gat426, gat407, gat408);
and 427gat (gat427, gat320, gat394, gat57);
assign gat428 = gat427;
assign gat429 = gat427;
assign gat430 = gat427;
assign gat431 = gat427;
and 432gat (gat432, gat395, gat24, gat288);
assign gat433 = gat432;
assign gat434 = gat432;
assign gat435 = gat432;
assign gat436 = gat432;
nand 437gat (gat437, gat396, gat289, gat58);
assign gat438 = gat437;
assign gat439 = gat437;
assign gat440 = gat437;
assign gat441 = gat437;
nand 442gat (gat442, gat375, gat67, gat158, gat397);
nand 443gat (gat443, gat398, gat321, gat25);
and 444gat (gat444, gat411, gat412);
and 445gat (gat445, gat414, gat415);
not 451gat (gat451, gat424);
assign gat452 = gat451;
assign gat453 = gat451;
assign gat454 = gat451;
assign gat455 = gat451;
assign gat456 = gat451;
assign gat457 = gat451;
assign gat458 = gat451;
assign gat459 = gat451;
nor 460gat (gat460, gat406, gat425);
assign gat461 = gat460;
assign gat462 = gat460;
nor 463gat (gat463, gat409, gat426);
assign gat464 = gat463;
assign gat465 = gat463;
nand 466gat (gat466, gat442, gat410);
assign gat467 = gat466;
assign gat468 = gat466;
assign gat469 = gat466;
assign gat470 = gat466;
assign gat471 = gat466;
assign gat472 = gat466;
assign gat473 = gat466;
assign gat474 = gat466;
and 475gat (gat475, gat144, gat428);
and 476gat (gat476, gat312, gat433);
and 477gat (gat477, gat147, gat429);
and 478gat (gat478, gat313, gat434);
and 479gat (gat479, gat150, gat430);
and 480gat (gat480, gat314, gat435);
and 481gat (gat481, gat154, gat431);
and 482gat (gat482, gat315, gat436);
nand 483gat (gat483, gat443, gat7);
assign gat484 = gat483;
assign gat485 = gat483;
assign gat486 = gat483;
assign gat487 = gat483;
or 488gat (gat488, gat371, gat438);
or 489gat (gat489, gat372, gat439);
or 490gat (gat490, gat373, gat440);
or 491gat (gat491, gat374, gat441);
nor 492gat (gat492, gat413, gat444);
assign gat493 = gat492;
assign gat494 = gat492;
nor 495gat (gat495, gat416, gat445);
assign gat496 = gat495;
assign gat497 = gat495;
nand 498gat (gat498, gat131, gat461);
or 499gat (gat499, gat132, gat462);
nand 500gat (gat500, gat464, gat136);
or 501gat (gat501, gat465, gat137);
and 502gat (gat502, gat95, gat467);
nor 503gat (gat503, gat475, gat476);
and 504gat (gat504, gat100, gat468);
nor 505gat (gat505, gat477, gat478);
and 506gat (gat506, gat105, gat469);
nor 507gat (gat507, gat479, gat480);
and 508gat (gat508, gat110, gat470);
nor 509gat (gat509, gat481, gat482);
and 510gat (gat510, gat145, gat484);
and 511gat (gat511, gat115, gat471);
and 512gat (gat512, gat148, gat485);
and 513gat (gat513, gat120, gat472);
and 514gat (gat514, gat151, gat486);
and 515gat (gat515, gat125, gat473);
and 516gat (gat516, gat155, gat487);
and 517gat (gat517, gat129, gat474);
nand 518gat (gat518, gat133, gat493);
or 519gat (gat519, gat134, gat494);
nand 520gat (gat520, gat496, gat208);
or 521gat (gat521, gat497, gat209);
and 522gat (gat522, gat452, gat162);
and 523gat (gat523, gat453, gat168);
and 524gat (gat524, gat454, gat174);
and 525gat (gat525, gat455, gat180);
and 526gat (gat526, gat456, gat186);
nand 527gat (gat527, gat457, gat192);
nand 528gat (gat528, gat458, gat198);
nand 529gat (gat529, gat459, gat204);
nand 530gat (gat530, gat498, gat499);
assign gat531 = gat530;
assign gat532 = gat530;
nand 533gat (gat533, gat500, gat501);
assign gat534 = gat533;
assign gat535 = gat533;
nor 536gat (gat536, gat309, gat502);
nor 537gat (gat537, gat316, gat504);
nor 538gat (gat538, gat317, gat506);
nor 539gat (gat539, gat318, gat508);
nor 540gat (gat540, gat510, gat511);
nor 541gat (gat541, gat512, gat513);
nor 542gat (gat542, gat514, gat515);
nor 543gat (gat543, gat516, gat517);
nand 544gat (gat544, gat518, gat519);
assign gat545 = gat544;
assign gat546 = gat544;
nand 547gat (gat547, gat520, gat521);
assign gat548 = gat547;
assign gat549 = gat547;
not 550gat (gat550, gat531);
not 551gat (gat551, gat534);
and 552gat (gat552, gat532, gat535);
nand 553gat (gat553, gat536, gat503);
assign gat554 = gat553;
assign gat555 = gat553;
assign gat556 = gat553;
nand 557gat (gat557, gat537, gat505);
assign gat558 = gat557;
assign gat559 = gat557;
assign gat560 = gat557;
nand 561gat (gat561, gat538, gat507);
assign gat562 = gat561;
assign gat563 = gat561;
assign gat564 = gat561;
nand 565gat (gat565, gat539, gat509);
assign gat566 = gat565;
assign gat567 = gat565;
assign gat568 = gat565;
nand 569gat (gat569, gat488, gat540);
assign gat570 = gat569;
assign gat571 = gat569;
assign gat572 = gat569;
nand 573gat (gat573, gat489, gat541);
assign gat574 = gat573;
assign gat575 = gat573;
assign gat576 = gat573;
nand 577gat (gat577, gat490, gat542);
assign gat578 = gat577;
assign gat579 = gat577;
assign gat580 = gat577;
nand 581gat (gat581, gat491, gat543);
assign gat582 = gat581;
assign gat583 = gat581;
assign gat584 = gat581;
not 585gat (gat585, gat545);
not 586gat (gat586, gat548);
and 587gat (gat587, gat546, gat549);
and 588gat (gat588, gat550, gat551);
and 589gat (gat589, gat585, gat586);
nand 590gat (gat590, gat554, gat163);
assign gat591 = gat590;
assign gat592 = gat590;
or 593gat (gat593, gat555, gat164);
assign gat594 = gat593;
assign gat595 = gat593;
and 596gat (gat596, gat247, gat556);
nand 597gat (gat597, gat558, gat169);
assign gat598 = gat597;
assign gat599 = gat597;
or 600gat (gat600, gat559, gat170);
assign gat601 = gat600;
assign gat602 = gat600;
assign gat603 = gat600;
assign gat604 = gat600;
and 605gat (gat605, gat248, gat560);
nand 606gat (gat606, gat562, gat175);
assign gat607 = gat606;
assign gat608 = gat606;
or 609gat (gat609, gat563, gat176);
assign gat610 = gat609;
assign gat611 = gat609;
assign gat612 = gat609;
assign gat613 = gat609;
assign gat614 = gat609;
and 615gat (gat615, gat249, gat564);
nand 616gat (gat616, gat566, gat181);
assign gat617 = gat616;
assign gat618 = gat616;
or 619gat (gat619, gat567, gat182);
assign gat620 = gat619;
assign gat621 = gat619;
assign gat622 = gat619;
assign gat623 = gat619;
and 624gat (gat624, gat250, gat568);
nand 625gat (gat625, gat570, gat187);
assign gat626 = gat625;
assign gat627 = gat625;
or 628gat (gat628, gat571, gat188);
assign gat629 = gat628;
assign gat630 = gat628;
and 631gat (gat631, gat251, gat572);
nand 632gat (gat632, gat574, gat193);
assign gat633 = gat632;
assign gat634 = gat632;
or 635gat (gat635, gat575, gat194);
assign gat636 = gat635;
assign gat637 = gat635;
assign gat638 = gat635;
assign gat639 = gat635;
and 640gat (gat640, gat252, gat576);
nand 641gat (gat641, gat578, gat199);
assign gat642 = gat641;
assign gat643 = gat641;
or 644gat (gat644, gat579, gat200);
assign gat645 = gat644;
assign gat646 = gat644;
assign gat647 = gat644;
assign gat648 = gat644;
assign gat649 = gat644;
and 650gat (gat650, gat253, gat580);
nand 651gat (gat651, gat582, gat205);
assign gat652 = gat651;
assign gat653 = gat651;
or 654gat (gat654, gat583, gat206);
assign gat655 = gat654;
assign gat656 = gat654;
assign gat657 = gat654;
assign gat658 = gat654;
and 659gat (gat659, gat254, gat584);
nor 660gat (gat660, gat552, gat588);
nor 661gat (gat661, gat587, gat589);
not 662gat (gat662, gat591);
assign gat663 = gat662;
assign gat664 = gat662;
and 665gat (gat665, gat594, gat592);
assign gat666 = gat665;
assign gat667 = gat665;
assign gat668 = gat665;
nor 669gat (gat669, gat596, gat522);
not 670gat (gat670, gat598);
assign gat671 = gat670;
assign gat672 = gat670;
and 673gat (gat673, gat601, gat599);
assign gat674 = gat673;
assign gat675 = gat673;
assign gat676 = gat673;
nor 677gat (gat677, gat605, gat523);
not 678gat (gat678, gat607);
assign gat679 = gat678;
assign gat680 = gat678;
assign gat681 = gat678;
and 682gat (gat682, gat610, gat608);
assign gat683 = gat682;
assign gat684 = gat682;
assign gat685 = gat682;
nor 686gat (gat686, gat615, gat524);
not 687gat (gat687, gat617);
assign gat688 = gat687;
assign gat689 = gat687;
assign gat690 = gat687;
assign gat691 = gat687;
and 692gat (gat692, gat620, gat618);
assign gat693 = gat692;
assign gat694 = gat692;
assign gat695 = gat692;
nor 696gat (gat696, gat624, gat525);
not 697gat (gat697, gat626);
assign gat698 = gat697;
assign gat699 = gat697;
and 700gat (gat700, gat629, gat627);
assign gat701 = gat700;
assign gat702 = gat700;
assign gat703 = gat700;
nor 704gat (gat704, gat631, gat526);
not 705gat (gat705, gat633);
assign gat706 = gat705;
assign gat707 = gat705;
and 708gat (gat708, gat636, gat634);
assign gat709 = gat708;
assign gat710 = gat708;
assign gat711 = gat708;
nor 712gat (gat712, gat337, gat640);
not 713gat (gat713, gat642);
assign gat714 = gat713;
assign gat715 = gat713;
assign gat716 = gat713;
and 717gat (gat717, gat645, gat643);
assign gat718 = gat717;
assign gat719 = gat717;
assign gat720 = gat717;
nor 721gat (gat721, gat339, gat650);
not 722gat (gat722, gat652);
assign gat723 = gat722;
assign gat724 = gat722;
assign gat725 = gat722;
assign gat726 = gat722;
and 727gat (gat727, gat655, gat653);
assign gat728 = gat727;
assign gat729 = gat727;
assign gat730 = gat727;
nor 731gat (gat731, gat341, gat659);
nand 732gat (gat732, gat656, gat262);
nand 733gat (gat733, gat646, gat657, gat263);
nand 734gat (gat734, gat637, gat647, gat658, gat264);
not 735gat (gat735, gat663);
and 736gat (gat736, gat229, gat666);
and 737gat (gat737, gat238, gat664);
not 738gat (gat738, gat671);
and 739gat (gat739, gat230, gat674);
and 740gat (gat740, gat239, gat672);
not 741gat (gat741, gat679);
and 742gat (gat742, gat231, gat683);
and 743gat (gat743, gat240, gat680);
not 744gat (gat744, gat688);
and 745gat (gat745, gat232, gat693);
and 746gat (gat746, gat241, gat689);
not 747gat (gat747, gat698);
and 748gat (gat748, gat233, gat701);
and 749gat (gat749, gat242, gat699);
not 750gat (gat750, gat706);
and 751gat (gat751, gat234, gat709);
and 752gat (gat752, gat243, gat707);
not 753gat (gat753, gat714);
and 754gat (gat754, gat235, gat718);
and 755gat (gat755, gat244, gat715);
not 756gat (gat756, gat723);
nor 757gat (gat757, gat728, gat265);
and 758gat (gat758, gat729, gat266);
and 759gat (gat759, gat236, gat730);
and 760gat (gat760, gat245, gat724);
nand 761gat (gat761, gat648, gat725);
nand 762gat (gat762, gat638, gat716);
nand 763gat (gat763, gat639, gat649, gat726);
nand 764gat (gat764, gat611, gat690);
nand 765gat (gat765, gat602, gat681);
nand 766gat (gat766, gat603, gat612, gat691);
nor 769gat (gat769, gat736, gat737);
nor 770gat (gat770, gat739, gat740);
nor 771gat (gat771, gat742, gat743);
nor 772gat (gat772, gat745, gat746);
nand 773gat (gat773, gat750, gat762, gat763, gat734);
assign gat774 = gat773;
assign gat775 = gat773;
assign gat776 = gat773;
nor 777gat (gat777, gat748, gat749);
nand 778gat (gat778, gat753, gat761, gat733);
assign gat779 = gat778;
assign gat780 = gat778;
nor 781gat (gat781, gat751, gat752);
nand 782gat (gat782, gat756, gat732);
assign gat783 = gat782;
assign gat784 = gat782;
nor 785gat (gat785, gat754, gat755);
nor 786gat (gat786, gat757, gat758);
nor 787gat (gat787, gat759, gat760);
nor 788gat (gat788, gat702, gat774);
and 789gat (gat789, gat703, gat775);
nor 790gat (gat790, gat710, gat779);
and 791gat (gat791, gat711, gat780);
nor 792gat (gat792, gat719, gat783);
and 793gat (gat793, gat720, gat784);
and 794gat (gat794, gat220, gat786);
nand 795gat (gat795, gat630, gat776);
nand 796gat (gat796, gat795, gat747);
assign gat797 = gat796;
assign gat798 = gat796;
assign gat799 = gat796;
assign gat800 = gat796;
assign gat801 = gat796;
nor 802gat (gat802, gat788, gat789);
nor 803gat (gat803, gat790, gat791);
nor 804gat (gat804, gat792, gat793);
nor 805gat (gat805, gat340, gat794);
nor 806gat (gat806, gat694, gat797);
and 807gat (gat807, gat695, gat798);
and 808gat (gat808, gat221, gat802);
and 809gat (gat809, gat222, gat803);
and 810gat (gat810, gat223, gat804);
nand 811gat (gat811, gat805, gat787, gat731, gat529);
nand 812gat (gat812, gat621, gat799);
nand 813gat (gat813, gat613, gat622, gat800);
nand 814gat (gat814, gat604, gat614, gat623, gat801);
nand 815gat (gat815, gat738, gat765, gat766, gat814);
assign gat816 = gat815;
assign gat817 = gat815;
assign gat818 = gat815;
nand 819gat (gat819, gat741, gat764, gat813);
assign gat820 = gat819;
assign gat821 = gat819;
nand 822gat (gat822, gat744, gat812);
assign gat823 = gat822;
assign gat824 = gat822;
nor 825gat (gat825, gat806, gat807);
nor 826gat (gat826, gat335, gat808);
nor 827gat (gat827, gat336, gat809);
nor 828gat (gat828, gat338, gat810);
not 829gat (gat829, gat811);
nor 830gat (gat830, gat667, gat816);
and 831gat (gat831, gat668, gat817);
nor 832gat (gat832, gat675, gat820);
and 833gat (gat833, gat676, gat821);
nor 834gat (gat834, gat684, gat823);
and 835gat (gat835, gat685, gat824);
and 836gat (gat836, gat224, gat825);
nand 837gat (gat837, gat826, gat777, gat704);
nand 838gat (gat838, gat827, gat781, gat712, gat527);
nand 839gat (gat839, gat828, gat785, gat721, gat528);
not 840gat (gat840, gat829);
nand 841gat (gat841, gat818, gat595);
nor 842gat (gat842, gat830, gat831);
nor 843gat (gat843, gat832, gat833);
nor 844gat (gat844, gat834, gat835);
nor 845gat (gat845, gat334, gat836);
not 846gat (gat846, gat837);
not 847gat (gat847, gat838);
not 848gat (gat848, gat839);
and 849gat (gat849, gat735, gat841);
and 851gat (gat851, gat225, gat842);
and 852gat (gat852, gat226, gat843);
and 853gat (gat853, gat227, gat844);
nand 854gat (gat854, gat845, gat772, gat696);
not 855gat (gat855, gat846);
not 856gat (gat856, gat847);
not 857gat (gat857, gat848);
not 858gat (gat858, gat849);
nor 859gat (gat859, gat417, gat851);
nor 860gat (gat860, gat332, gat852);
nor 861gat (gat861, gat333, gat853);
not 862gat (gat862, gat854);
nand 867gat (gat867, gat859, gat769, gat669);
nand 868gat (gat868, gat860, gat770, gat677);
nand 869gat (gat869, gat861, gat771, gat686);
not 870gat (gat870, gat862);
not 871gat (gat871, gat867);
not 872gat (gat872, gat868);
not 873gat (gat873, gat869);
not 875gat (gat875, gat871);
not 876gat (gat876, gat872);
not 877gat (gat877, gat873);
endmodule